.include sqj960ep_ps.txt


.SUBCKT SQJ476ELP D1 G1 S1 D2 G2 S2
X1 D1 G1 S1 SQJ960EP
X2 D2 G2 S2 SQJ960EP
.ENDS
